// модуль, который реализует расширенение
// 16-битной знаковой константы до 32-битной
module sign_extend(in, out);
  input [15:0] in;
  output [31:0] out;

  //assign out = {{16{in[15]}}, in};
  assign out[15:0] = in;
  assign out[16] = in[15] == 1;
  assign out[17] = in[15] == 1;
  assign out[18] = in[15] == 1;
  assign out[19] = in[15] == 1;
  assign out[20] = in[15] == 1;
  assign out[21] = in[15] == 1;
  assign out[22] = in[15] == 1;
  assign out[23] = in[15] == 1;
  assign out[24] = in[15] == 1;
  assign out[25] = in[15] == 1;
  assign out[26] = in[15] == 1;
  assign out[27] = in[15] == 1;
  assign out[28] = in[15] == 1;
  assign out[29] = in[15] == 1;
  assign out[30] = in[15] == 1;
  assign out[31] = in[15] == 1;
endmodule

// модуль, который реализует побитовый сдвиг числа
// влево на 2 бита
module shl_2(in, out);
  input [31:0] in;
  output [31:0] out;

  assign out[31:2] = in[29:0];
  assign out[1:0] = 2'b00;
endmodule

// 32 битный сумматор
module adder(a, b, out);
  input [31:0] a, b;
  output [31:0] out;

  assign out = a + b;
endmodule

// 32-битный мультиплексор
module mux2_32(d0, d1, a, out);
  input [31:0] d0, d1;
  input a;
  output [31:0] out;
  assign out = a ? d1 : d0;
endmodule

// 5 - битный мультиплексор
module mux2_5(d0, d1, a, out);
  input [4:0] d0, d1;
  input a;
  output [4:0] out;
  assign out = a ? d1 : d0;
endmodule

module and_gate(a, b, out);
  input wire a, b;
  output wire out;

  wire nand_out;

  nand_gate nand_gate1(a, b, nand_out);
  not_gate not_gate1(nand_out, out);
endmodule

module nand_gate(a, b, out);
  input wire a, b;
  output out;

  supply1 pwr;
  supply0 gnd;

  wire nmos1_out;

  pmos pmos1(out, pwr, a);
  pmos pmos2(out, pwr, b);

  nmos nmos1(nmos1_out, gnd, b);
  nmos nmos2(out, nmos1_out, a);
  // pmos pmos1(out, pwr, a);
  // nmos nmos1(out, gnd, a);
endmodule


module not_gate(a, out);
  input wire a;
  output out;

  supply1 pwr;
  supply0 gnd;

  // 1 - сток, 2 - исток, 3 - база
  pmos pmos1(out, pwr, a);
  nmos nmos1(out, gnd, a);
endmodule

module or_gate(a, b, out);
  input a, b;
  output out;

  wire na, nb;

  not_gate nt1(a, na);
  not_gate nt2(b, nb);

  nand_gate nand1(na, nb, out);
endmodule

